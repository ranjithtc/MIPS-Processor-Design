library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity imem is
    Port ( a : in  STD_LOGIC_VECTOR (5 downto 0);
           rd : out  STD_LOGIC_VECTOR (31 downto 0));
end imem;

architecture Behavioral of imem is
	type mem is array(0 to 63) of std_logic_vector(31 downto 0);
	constant code : mem:=(

		-- Load here your software.
		
x"20020005", -- 001000 00000000100000000000000101
x"2003000c", -- 001000 00000000110000000000001100
x"2067fff7", -- 001000 00011001111111111111110111
x"00e22025", -- 000000 00111000100010000000100101
x"00642824", -- 000000 00011001000010100000100100
x"00a42820", -- 000000 00101001000010100000100000
x"10a7000a", -- 000100 00101001110000000000001010  -- beq
x"0064202a", -- 000000 00011001000010000000101010 
x"10800001", -- 000100 00100000000000000000000001  -- beq
x"20050000", -- 001000 00000001010000000000000000  -- shouldnt happen because branch taken 
x"00e2202a", -- 000000 00111000100010000000101010  
x"00853820", -- 000000 00100001010011100000100000
x"00e23822", -- 000000 00111000100011100000100010
x"ac670044", -- 101011 00011001110000000001000100
x"8c020050", -- 100011 00000000100000000001010000
x"08000011", -- 000010 00000000000000000000010001  -- j
x"20020001", -- 001000 00000000100000000000000001  -- shouldnt happen because of jump
x"ac020054", -- 101011 00000000100000000001010100

	others=> x"00000000");

begin

rd <= code(to_integer(unsigned(a)));

end Behavioral;